`timescale 1ns / 1ps

module mult(
	input mul_clk,
	input resetn,
	input mul_signed,
	input [31:0] x,
	input [31:0] y,

	output [63:0] result
);
  wire [63:0] p00, p01, p02, p03, p04, p05, p06, p07, p08;
  wire [63:0] p09, p10, p11, p12, p13, p14, p15, p16;
  wire        c00, c01, c02, c03, c04, c05, c06, c07, c08;
  wire        c09, c10, c11, c12, c13, c14, c15, c16;
  
  wire [16:0] N00, N01, N02, N03, N04, N05, N06, N07;
  wire [16:0] N08, N09, N10, N11, N12, N13, N14, N15;
  wire [16:0] N16, N17, N18, N19, N20, N21, N22, N23;
  wire [16:0] N24, N25, N26, N27, N28, N29, N30, N31;
  wire [16:0] N32, N33, N34, N35, N36, N37, N38, N39;
  wire [16:0] N40, N41, N42, N43, N44, N45, N46, N47;
  wire [16:0] N48, N49, N50, N51, N52, N53, N54, N55;
  wire [16:0] N56, N57, N58, N59, N60, N61, N62, N63;
  wire [16:0] C;

  wire [63:0] C_wallace;
  wire [63:0] S_wallace;
  
  reg  [63:0] final_S;
  reg  [63:0] final_C;
  reg         final_Cin;
  wire [63:0] final_result;
  
  wire [33:0] A;
  wire [33:0] B; 
  
  assign A = (mul_signed)? {{2{x[31]}}, x} : {2'b00, x};
  assign B = (mul_signed)? {{2{y[31]}}, y} : {2'b00, y};
  
  assign result = final_result;
	always@(posedge mul_clk)
	begin
	  if(!resetn) begin
	    final_S   <= 64'b0;
	    final_C   <= 64'b0;
	    final_Cin <=  1'b0;
	  end
	  else begin
	    final_S   <= S_wallace;
	    final_C   <= {C_wallace[62:0],C[14]};
	    final_Cin <= C[15];
	  end
	end

  assign C = {c16, c15, c14, c13, c12, c11, c10, c09, c08, c07, c06, c05, c04, c03, c02, c01, c00};
  
  booth booth(.A(A), .B(B),
              .p00(p00), .p01(p01), .p02(p02), .p03(p03), .p04(p04), .p05(p05), .p06(p06), .p07(p07), .p08(p08),
              .p09(p09), .p10(p10), .p11(p11), .p12(p12), .p13(p13), .p14(p14), .p15(p15), .p16(p16), 
              .c00(c00), .c01(c01), .c02(c02), .c03(c03), .c04(c04), .c05(c05), .c06(c06), .c07(c07), .c08(c08),
              .c09(c09), .c10(c10), .c11(c11), .c12(c12), .c13(c13), .c14(c14), .c15(c15), .c16(c16)
              );

  switch switch(
              .p00(p00), .p01(p01), .p02(p02), .p03(p03), .p04(p04), .p05(p05), .p06(p06), .p07(p07), .p08(p08),
              .p09(p09), .p10(p10), .p11(p11), .p12(p12), .p13(p13), .p14(p14), .p15(p15), .p16(p16),
              
              .N00(N00), .N01(N01), .N02(N02), .N03(N03), .N04(N04), .N05(N05), .N06(N06), .N07(N07), 
              .N08(N08), .N09(N09), .N10(N10), .N11(N11), .N12(N12), .N13(N13), .N14(N14), .N15(N15), 
              .N16(N16), .N17(N17), .N18(N18), .N19(N19), .N20(N20), .N21(N21), .N22(N22), .N23(N23),
              .N24(N24), .N25(N25), .N26(N26), .N27(N27), .N28(N28), .N29(N29), .N30(N30), .N31(N31), 
              .N32(N32), .N33(N33), .N34(N34), .N35(N35), .N36(N36), .N37(N37), .N38(N38), .N39(N39), 
              .N40(N40), .N41(N41), .N42(N42), .N43(N43), .N44(N44), .N45(N45), .N46(N46), .N47(N47), 
              .N48(N48), .N49(N49), .N50(N50), .N51(N51), .N52(N52), .N53(N53), .N54(N54), .N55(N55), 
              .N56(N56), .N57(N57), .N58(N58), .N59(N59), .N60(N60), .N61(N61), .N62(N62), .N63(N63)
              );
              
  Wallace Wallace(
              .N00(N00), .N01(N01), .N02(N02), .N03(N03), .N04(N04), .N05(N05), .N06(N06), .N07(N07), 
              .N08(N08), .N09(N09), .N10(N10), .N11(N11), .N12(N12), .N13(N13), .N14(N14), .N15(N15), 
              .N16(N16), .N17(N17), .N18(N18), .N19(N19), .N20(N20), .N21(N21), .N22(N22), .N23(N23),
              .N24(N24), .N25(N25), .N26(N26), .N27(N27), .N28(N28), .N29(N29), .N30(N30), .N31(N31), 
              .N32(N32), .N33(N33), .N34(N34), .N35(N35), .N36(N36), .N37(N37), .N38(N38), .N39(N39), 
              .N40(N40), .N41(N41), .N42(N42), .N43(N43), .N44(N44), .N45(N45), .N46(N46), .N47(N47), 
              .N48(N48), .N49(N49), .N50(N50), .N51(N51), .N52(N52), .N53(N53), .N54(N54), .N55(N55), 
              .N56(N56), .N57(N57), .N58(N58), .N59(N59), .N60(N60), .N61(N61), .N62(N62), .N63(N63),
              .Cin(C[13:0]),

              .Cout(C_wallace),
              .S(S_wallace)
              );
             
  final_adder adder(.A(final_S), .B(final_C), .Cin(final_Cin), .result(final_result));
endmodule



module booth(
  input  [33:0] A,
  input  [33:0] B,

  output [63:0] p00, p01, p02, p03, p04, p05, p06, p07, p08,
  output [63:0] p09, p10, p11, p12, p13, p14, p15, p16,
  output        c00, c01, c02, c03, c04, c05, c06, c07, c08,
  output        c09, c10, c11, c12, c13, c14, c15, c16
  
);

  partial_product p_prod00(.A(A), .B({B[ 1: 0],1'b0}), .shift(6'd00), .p(p00), .c(c00)),
                  p_prod01(.A(A), .B( B[ 3: 1]      ), .shift(6'd02), .p(p01), .c(c01)),
                  p_prod02(.A(A), .B( B[ 5: 3]      ), .shift(6'd04), .p(p02), .c(c02)),
                  p_prod03(.A(A), .B( B[ 7: 5]      ), .shift(6'd06), .p(p03), .c(c03)),
                  p_prod04(.A(A), .B( B[ 9: 7]      ), .shift(6'd08), .p(p04), .c(c04)),
                  p_prod05(.A(A), .B( B[11: 9]      ), .shift(6'd10), .p(p05), .c(c05)),
                  p_prod06(.A(A), .B( B[13:11]      ), .shift(6'd12), .p(p06), .c(c06)),
                  p_prod07(.A(A), .B( B[15:13]      ), .shift(6'd14), .p(p07), .c(c07)),
                  p_prod08(.A(A), .B( B[17:15]      ), .shift(6'd16), .p(p08), .c(c08)),
                  p_prod09(.A(A), .B( B[19:17]      ), .shift(6'd18), .p(p09), .c(c09)),
                  p_prod10(.A(A), .B( B[21:19]      ), .shift(6'd20), .p(p10), .c(c10)),
                  p_prod11(.A(A), .B( B[23:21]      ), .shift(6'd22), .p(p11), .c(c11)),
                  p_prod12(.A(A), .B( B[25:23]      ), .shift(6'd24), .p(p12), .c(c12)),
                  p_prod13(.A(A), .B( B[27:25]      ), .shift(6'd26), .p(p13), .c(c13)),
                  p_prod14(.A(A), .B( B[29:27]      ), .shift(6'd28), .p(p14), .c(c14)),
                  p_prod15(.A(A), .B( B[31:29]      ), .shift(6'd30), .p(p15), .c(c15)),
                  p_prod16(.A(A), .B( B[33:31]      ), .shift(6'd32), .p(p16), .c(c16));
endmodule
 
module partial_product(
  input  [33:0] A,
  input  [ 2:0] B,
  input  [ 5:0] shift,
  
  output [63:0] p,
  output        c
);

  wire [33:0] p_temp;
  wire [95:0] p_pre;
  wire [33:0] A_neg;
  
  assign A_neg = ~A;

  assign p_temp = (B==3'b001)? A:
                  (B==3'b010)? A:
                  (B==3'b011)? {A[32:0], 1'b0}:
                  (B==3'b100)? {A_neg[32:0], 1'b1}:
                  (B==3'b101)? A_neg:
                  (B==3'b110)? A_neg:
                               34'b0;
                               
  assign c = (B==3'b100||B==3'b101||B==3'b110)? 1'b1 : 1'b0;
  
  assign p_pre = {{30{p_temp[33]}}, p_temp, {32{c}}} << shift;

  assign p = p_pre[95:32];                

endmodule


module switch(
  input  [63:0] p00, p01, p02, p03, p04, p05, p06, p07, p08,
  input  [63:0] p09, p10, p11, p12, p13, p14, p15, p16,
  
  output [16:0] N00, N01, N02, N03, N04, N05, N06, N07,
  output [16:0] N08, N09, N10, N11, N12, N13, N14, N15,
  output [16:0] N16, N17, N18, N19, N20, N21, N22, N23,
  output [16:0] N24, N25, N26, N27, N28, N29, N30, N31,
  output [16:0] N32, N33, N34, N35, N36, N37, N38, N39,
  output [16:0] N40, N41, N42, N43, N44, N45, N46, N47,
  output [16:0] N48, N49, N50, N51, N52, N53, N54, N55,
  output [16:0] N56, N57, N58, N59, N60, N61, N62, N63
);

  assign N00 = {p00[00], p01[00] ,p02[00], p03[00], p04[00], p05[00], p06[00], p07[00], p08[00], p09[00], p10[00], p11[00], p12[00], p13[00], p14[00], p15[00], p16[00]};
  assign N01 = {p00[01], p01[01] ,p02[01], p03[01], p04[01], p05[01], p06[01], p07[01], p08[01], p09[01], p10[01], p11[01], p12[01], p13[01], p14[01], p15[01], p16[01]};
  assign N02 = {p00[02], p01[02] ,p02[02], p03[02], p04[02], p05[02], p06[02], p07[02], p08[02], p09[02], p10[02], p11[02], p12[02], p13[02], p14[02], p15[02], p16[02]};
  assign N03 = {p00[03], p01[03] ,p02[03], p03[03], p04[03], p05[03], p06[03], p07[03], p08[03], p09[03], p10[03], p11[03], p12[03], p13[03], p14[03], p15[03], p16[03]};
  assign N04 = {p00[04], p01[04] ,p02[04], p03[04], p04[04], p05[04], p06[04], p07[04], p08[04], p09[04], p10[04], p11[04], p12[04], p13[04], p14[04], p15[04], p16[04]};
  assign N05 = {p00[05], p01[05] ,p02[05], p03[05], p04[05], p05[05], p06[05], p07[05], p08[05], p09[05], p10[05], p11[05], p12[05], p13[05], p14[05], p15[05], p16[05]};
  assign N06 = {p00[06], p01[06] ,p02[06], p03[06], p04[06], p05[06], p06[06], p07[06], p08[06], p09[06], p10[06], p11[06], p12[06], p13[06], p14[06], p15[06], p16[06]};
  assign N07 = {p00[07], p01[07] ,p02[07], p03[07], p04[07], p05[07], p06[07], p07[07], p08[07], p09[07], p10[07], p11[07], p12[07], p13[07], p14[07], p15[07], p16[07]};
  assign N08 = {p00[08], p01[08] ,p02[08], p03[08], p04[08], p05[08], p06[08], p07[08], p08[08], p09[08], p10[08], p11[08], p12[08], p13[08], p14[08], p15[08], p16[08]};
  assign N09 = {p00[09], p01[09] ,p02[09], p03[09], p04[09], p05[09], p06[09], p07[09], p08[09], p09[09], p10[09], p11[09], p12[09], p13[09], p14[09], p15[09], p16[09]};
  assign N10 = {p00[10], p01[10] ,p02[10], p03[10], p04[10], p05[10], p06[10], p07[10], p08[10], p09[10], p10[10], p11[10], p12[10], p13[10], p14[10], p15[10], p16[10]};
  assign N11 = {p00[11], p01[11] ,p02[11], p03[11], p04[11], p05[11], p06[11], p07[11], p08[11], p09[11], p10[11], p11[11], p12[11], p13[11], p14[11], p15[11], p16[11]};
  assign N12 = {p00[12], p01[12] ,p02[12], p03[12], p04[12], p05[12], p06[12], p07[12], p08[12], p09[12], p10[12], p11[12], p12[12], p13[12], p14[12], p15[12], p16[12]};
  assign N13 = {p00[13], p01[13] ,p02[13], p03[13], p04[13], p05[13], p06[13], p07[13], p08[13], p09[13], p10[13], p11[13], p12[13], p13[13], p14[13], p15[13], p16[13]};
  assign N14 = {p00[14], p01[14] ,p02[14], p03[14], p04[14], p05[14], p06[14], p07[14], p08[14], p09[14], p10[14], p11[14], p12[14], p13[14], p14[14], p15[14], p16[14]};
  assign N15 = {p00[15], p01[15] ,p02[15], p03[15], p04[15], p05[15], p06[15], p07[15], p08[15], p09[15], p10[15], p11[15], p12[15], p13[15], p14[15], p15[15], p16[15]};
  assign N16 = {p00[16], p01[16] ,p02[16], p03[16], p04[16], p05[16], p06[16], p07[16], p08[16], p09[16], p10[16], p11[16], p12[16], p13[16], p14[16], p15[16], p16[16]};
  assign N17 = {p00[17], p01[17] ,p02[17], p03[17], p04[17], p05[17], p06[17], p07[17], p08[17], p09[17], p10[17], p11[17], p12[17], p13[17], p14[17], p15[17], p16[17]};
  assign N18 = {p00[18], p01[18] ,p02[18], p03[18], p04[18], p05[18], p06[18], p07[18], p08[18], p09[18], p10[18], p11[18], p12[18], p13[18], p14[18], p15[18], p16[18]};
  assign N19 = {p00[19], p01[19] ,p02[19], p03[19], p04[19], p05[19], p06[19], p07[19], p08[19], p09[19], p10[19], p11[19], p12[19], p13[19], p14[19], p15[19], p16[19]};
  assign N20 = {p00[20], p01[20] ,p02[20], p03[20], p04[20], p05[20], p06[20], p07[20], p08[20], p09[20], p10[20], p11[20], p12[20], p13[20], p14[20], p15[20], p16[20]};
  assign N21 = {p00[21], p01[21] ,p02[21], p03[21], p04[21], p05[21], p06[21], p07[21], p08[21], p09[21], p10[21], p11[21], p12[21], p13[21], p14[21], p15[21], p16[21]};
  assign N22 = {p00[22], p01[22] ,p02[22], p03[22], p04[22], p05[22], p06[22], p07[22], p08[22], p09[22], p10[22], p11[22], p12[22], p13[22], p14[22], p15[22], p16[22]};
  assign N23 = {p00[23], p01[23] ,p02[23], p03[23], p04[23], p05[23], p06[23], p07[23], p08[23], p09[23], p10[23], p11[23], p12[23], p13[23], p14[23], p15[23], p16[23]};
  assign N24 = {p00[24], p01[24] ,p02[24], p03[24], p04[24], p05[24], p06[24], p07[24], p08[24], p09[24], p10[24], p11[24], p12[24], p13[24], p14[24], p15[24], p16[24]};
  assign N25 = {p00[25], p01[25] ,p02[25], p03[25], p04[25], p05[25], p06[25], p07[25], p08[25], p09[25], p10[25], p11[25], p12[25], p13[25], p14[25], p15[25], p16[25]};
  assign N26 = {p00[26], p01[26] ,p02[26], p03[26], p04[26], p05[26], p06[26], p07[26], p08[26], p09[26], p10[26], p11[26], p12[26], p13[26], p14[26], p15[26], p16[26]};
  assign N27 = {p00[27], p01[27] ,p02[27], p03[27], p04[27], p05[27], p06[27], p07[27], p08[27], p09[27], p10[27], p11[27], p12[27], p13[27], p14[27], p15[27], p16[27]};
  assign N28 = {p00[28], p01[28] ,p02[28], p03[28], p04[28], p05[28], p06[28], p07[28], p08[28], p09[28], p10[28], p11[28], p12[28], p13[28], p14[28], p15[28], p16[28]};
  assign N29 = {p00[29], p01[29] ,p02[29], p03[29], p04[29], p05[29], p06[29], p07[29], p08[29], p09[29], p10[29], p11[29], p12[29], p13[29], p14[29], p15[29], p16[29]};
  assign N30 = {p00[30], p01[30] ,p02[30], p03[30], p04[30], p05[30], p06[30], p07[30], p08[30], p09[30], p10[30], p11[30], p12[30], p13[30], p14[30], p15[30], p16[30]};
  assign N31 = {p00[31], p01[31] ,p02[31], p03[31], p04[31], p05[31], p06[31], p07[31], p08[31], p09[31], p10[31], p11[31], p12[31], p13[31], p14[31], p15[31], p16[31]};
  assign N32 = {p00[32], p01[32] ,p02[32], p03[32], p04[32], p05[32], p06[32], p07[32], p08[32], p09[32], p10[32], p11[32], p12[32], p13[32], p14[32], p15[32], p16[32]};
  assign N33 = {p00[33], p01[33] ,p02[33], p03[33], p04[33], p05[33], p06[33], p07[33], p08[33], p09[33], p10[33], p11[33], p12[33], p13[33], p14[33], p15[33], p16[33]};
  assign N34 = {p00[34], p01[34] ,p02[34], p03[34], p04[34], p05[34], p06[34], p07[34], p08[34], p09[34], p10[34], p11[34], p12[34], p13[34], p14[34], p15[34], p16[34]};
  assign N35 = {p00[35], p01[35] ,p02[35], p03[35], p04[35], p05[35], p06[35], p07[35], p08[35], p09[35], p10[35], p11[35], p12[35], p13[35], p14[35], p15[35], p16[35]};
  assign N36 = {p00[36], p01[36] ,p02[36], p03[36], p04[36], p05[36], p06[36], p07[36], p08[36], p09[36], p10[36], p11[36], p12[36], p13[36], p14[36], p15[36], p16[36]};
  assign N37 = {p00[37], p01[37] ,p02[37], p03[37], p04[37], p05[37], p06[37], p07[37], p08[37], p09[37], p10[37], p11[37], p12[37], p13[37], p14[37], p15[37], p16[37]};
  assign N38 = {p00[38], p01[38] ,p02[38], p03[38], p04[38], p05[38], p06[38], p07[38], p08[38], p09[38], p10[38], p11[38], p12[38], p13[38], p14[38], p15[38], p16[38]};
  assign N39 = {p00[39], p01[39] ,p02[39], p03[39], p04[39], p05[39], p06[39], p07[39], p08[39], p09[39], p10[39], p11[39], p12[39], p13[39], p14[39], p15[39], p16[39]};
  assign N40 = {p00[40], p01[40] ,p02[40], p03[40], p04[40], p05[40], p06[40], p07[40], p08[40], p09[40], p10[40], p11[40], p12[40], p13[40], p14[40], p15[40], p16[40]};
  assign N41 = {p00[41], p01[41] ,p02[41], p03[41], p04[41], p05[41], p06[41], p07[41], p08[41], p09[41], p10[41], p11[41], p12[41], p13[41], p14[41], p15[41], p16[41]};
  assign N42 = {p00[42], p01[42] ,p02[42], p03[42], p04[42], p05[42], p06[42], p07[42], p08[42], p09[42], p10[42], p11[42], p12[42], p13[42], p14[42], p15[42], p16[42]};
  assign N43 = {p00[43], p01[43] ,p02[43], p03[43], p04[43], p05[43], p06[43], p07[43], p08[43], p09[43], p10[43], p11[43], p12[43], p13[43], p14[43], p15[43], p16[43]};
  assign N44 = {p00[44], p01[44] ,p02[44], p03[44], p04[44], p05[44], p06[44], p07[44], p08[44], p09[44], p10[44], p11[44], p12[44], p13[44], p14[44], p15[44], p16[44]};
  assign N45 = {p00[45], p01[45] ,p02[45], p03[45], p04[45], p05[45], p06[45], p07[45], p08[45], p09[45], p10[45], p11[45], p12[45], p13[45], p14[45], p15[45], p16[45]};
  assign N46 = {p00[46], p01[46] ,p02[46], p03[46], p04[46], p05[46], p06[46], p07[46], p08[46], p09[46], p10[46], p11[46], p12[46], p13[46], p14[46], p15[46], p16[46]};
  assign N47 = {p00[47], p01[47] ,p02[47], p03[47], p04[47], p05[47], p06[47], p07[47], p08[47], p09[47], p10[47], p11[47], p12[47], p13[47], p14[47], p15[47], p16[47]};
  assign N48 = {p00[48], p01[48] ,p02[48], p03[48], p04[48], p05[48], p06[48], p07[48], p08[48], p09[48], p10[48], p11[48], p12[48], p13[48], p14[48], p15[48], p16[48]};
  assign N49 = {p00[49], p01[49] ,p02[49], p03[49], p04[49], p05[49], p06[49], p07[49], p08[49], p09[49], p10[49], p11[49], p12[49], p13[49], p14[49], p15[49], p16[49]};
  assign N50 = {p00[50], p01[50] ,p02[50], p03[50], p04[50], p05[50], p06[50], p07[50], p08[50], p09[50], p10[50], p11[50], p12[50], p13[50], p14[50], p15[50], p16[50]};
  assign N51 = {p00[51], p01[51] ,p02[51], p03[51], p04[51], p05[51], p06[51], p07[51], p08[51], p09[51], p10[51], p11[51], p12[51], p13[51], p14[51], p15[51], p16[51]};
  assign N52 = {p00[52], p01[52] ,p02[52], p03[52], p04[52], p05[52], p06[52], p07[52], p08[52], p09[52], p10[52], p11[52], p12[52], p13[52], p14[52], p15[52], p16[52]};
  assign N53 = {p00[53], p01[53] ,p02[53], p03[53], p04[53], p05[53], p06[53], p07[53], p08[53], p09[53], p10[53], p11[53], p12[53], p13[53], p14[53], p15[53], p16[53]};
  assign N54 = {p00[54], p01[54] ,p02[54], p03[54], p04[54], p05[54], p06[54], p07[54], p08[54], p09[54], p10[54], p11[54], p12[54], p13[54], p14[54], p15[54], p16[54]};
  assign N55 = {p00[55], p01[55] ,p02[55], p03[55], p04[55], p05[55], p06[55], p07[55], p08[55], p09[55], p10[55], p11[55], p12[55], p13[55], p14[55], p15[55], p16[55]};
  assign N56 = {p00[56], p01[56] ,p02[56], p03[56], p04[56], p05[56], p06[56], p07[56], p08[56], p09[56], p10[56], p11[56], p12[56], p13[56], p14[56], p15[56], p16[56]};
  assign N57 = {p00[57], p01[57] ,p02[57], p03[57], p04[57], p05[57], p06[57], p07[57], p08[57], p09[57], p10[57], p11[57], p12[57], p13[57], p14[57], p15[57], p16[57]};
  assign N58 = {p00[58], p01[58] ,p02[58], p03[58], p04[58], p05[58], p06[58], p07[58], p08[58], p09[58], p10[58], p11[58], p12[58], p13[58], p14[58], p15[58], p16[58]};
  assign N59 = {p00[59], p01[59] ,p02[59], p03[59], p04[59], p05[59], p06[59], p07[59], p08[59], p09[59], p10[59], p11[59], p12[59], p13[59], p14[59], p15[59], p16[59]};
  assign N60 = {p00[60], p01[60] ,p02[60], p03[60], p04[60], p05[60], p06[60], p07[60], p08[60], p09[60], p10[60], p11[60], p12[60], p13[60], p14[60], p15[60], p16[60]};
  assign N61 = {p00[61], p01[61] ,p02[61], p03[61], p04[61], p05[61], p06[61], p07[61], p08[61], p09[61], p10[61], p11[61], p12[61], p13[61], p14[61], p15[61], p16[61]};
  assign N62 = {p00[62], p01[62] ,p02[62], p03[62], p04[62], p05[62], p06[62], p07[62], p08[62], p09[62], p10[62], p11[62], p12[62], p13[62], p14[62], p15[62], p16[62]};
  assign N63 = {p00[63], p01[63] ,p02[63], p03[63], p04[63], p05[63], p06[63], p07[63], p08[63], p09[63], p10[63], p11[63], p12[63], p13[63], p14[63], p15[63], p16[63]};

endmodule 

module Wallace (
  input  [16:0] N00, N01, N02, N03, N04, N05, N06, N07,
  input  [16:0] N08, N09, N10, N11, N12, N13, N14, N15,
  input  [16:0] N16, N17, N18, N19, N20, N21, N22, N23,
  input  [16:0] N24, N25, N26, N27, N28, N29, N30, N31,
  input  [16:0] N32, N33, N34, N35, N36, N37, N38, N39,
  input  [16:0] N40, N41, N42, N43, N44, N45, N46, N47,
  input  [16:0] N48, N49, N50, N51, N52, N53, N54, N55,
  input  [16:0] N56, N57, N58, N59, N60, N61, N62, N63,
  input  [13:0] Cin,

  output [63:0] Cout,
  output [63:0] S
  );
  
  wire [13:0] Cout00, Cout01, Cout02, Cout03, Cout04, Cout05, Cout06, Cout07, Cout08, Cout09;
  wire [13:0] Cout10, Cout11, Cout12, Cout13, Cout14, Cout15, Cout16, Cout17, Cout18, Cout19;
  wire [13:0] Cout20, Cout21, Cout22, Cout23, Cout24, Cout25, Cout26, Cout27, Cout28, Cout29;
  wire [13:0] Cout30, Cout31, Cout32, Cout33, Cout34, Cout35, Cout36, Cout37, Cout38, Cout39;
  wire [13:0] Cout40, Cout41, Cout42, Cout43, Cout44, Cout45, Cout46, Cout47, Cout48, Cout49;
  wire [13:0] Cout50, Cout51, Cout52, Cout53, Cout54, Cout55, Cout56, Cout57, Cout58, Cout59;
  wire [13:0] Cout60, Cout61, Cout62, Cout63;
  
  
  one_bit_Wallace_tree tree00(.N(N00), .Cin(Cin    ), .Cout(Cout00), .C(Cout[00]), .S(S[00])),
                       tree01(.N(N01), .Cin(Cout00 ), .Cout(Cout01), .C(Cout[01]), .S(S[01])),
                       tree02(.N(N02), .Cin(Cout01 ), .Cout(Cout02), .C(Cout[02]), .S(S[02])),
                       tree03(.N(N03), .Cin(Cout02 ), .Cout(Cout03), .C(Cout[03]), .S(S[03])),
                       tree04(.N(N04), .Cin(Cout03 ), .Cout(Cout04), .C(Cout[04]), .S(S[04])),
                       tree05(.N(N05), .Cin(Cout04 ), .Cout(Cout05), .C(Cout[05]), .S(S[05])),
                       tree06(.N(N06), .Cin(Cout05 ), .Cout(Cout06), .C(Cout[06]), .S(S[06])),
                       tree07(.N(N07), .Cin(Cout06 ), .Cout(Cout07), .C(Cout[07]), .S(S[07])),
                       tree08(.N(N08), .Cin(Cout07 ), .Cout(Cout08), .C(Cout[08]), .S(S[08])),
                       tree09(.N(N09), .Cin(Cout08 ), .Cout(Cout09), .C(Cout[09]), .S(S[09])),
                       
                       tree10(.N(N10), .Cin(Cout09 ), .Cout(Cout10), .C(Cout[10]), .S(S[10])),
                       tree11(.N(N11), .Cin(Cout10 ), .Cout(Cout11), .C(Cout[11]), .S(S[11])),
                       tree12(.N(N12), .Cin(Cout11 ), .Cout(Cout12), .C(Cout[12]), .S(S[12])),
                       tree13(.N(N13), .Cin(Cout12 ), .Cout(Cout13), .C(Cout[13]), .S(S[13])),
                       tree14(.N(N14), .Cin(Cout13 ), .Cout(Cout14), .C(Cout[14]), .S(S[14])),
                       tree15(.N(N15), .Cin(Cout14 ), .Cout(Cout15), .C(Cout[15]), .S(S[15])),
                       tree16(.N(N16), .Cin(Cout15 ), .Cout(Cout16), .C(Cout[16]), .S(S[16])),
                       tree17(.N(N17), .Cin(Cout16 ), .Cout(Cout17), .C(Cout[17]), .S(S[17])),
                       tree18(.N(N18), .Cin(Cout17 ), .Cout(Cout18), .C(Cout[18]), .S(S[18])),
                       tree19(.N(N19), .Cin(Cout18 ), .Cout(Cout19), .C(Cout[19]), .S(S[19])),
                       
                       tree20(.N(N20), .Cin(Cout19 ), .Cout(Cout20), .C(Cout[20]), .S(S[20])),
                       tree21(.N(N21), .Cin(Cout20 ), .Cout(Cout21), .C(Cout[21]), .S(S[21])),
                       tree22(.N(N22), .Cin(Cout21 ), .Cout(Cout22), .C(Cout[22]), .S(S[22])),
                       tree23(.N(N23), .Cin(Cout22 ), .Cout(Cout23), .C(Cout[23]), .S(S[23])),
                       tree24(.N(N24), .Cin(Cout23 ), .Cout(Cout24), .C(Cout[24]), .S(S[24])),
                       tree25(.N(N25), .Cin(Cout24 ), .Cout(Cout25), .C(Cout[25]), .S(S[25])),
                       tree26(.N(N26), .Cin(Cout25 ), .Cout(Cout26), .C(Cout[26]), .S(S[26])),
                       tree27(.N(N27), .Cin(Cout26 ), .Cout(Cout27), .C(Cout[27]), .S(S[27])),
                       tree28(.N(N28), .Cin(Cout27 ), .Cout(Cout28), .C(Cout[28]), .S(S[28])),
                       tree29(.N(N29), .Cin(Cout28 ), .Cout(Cout29), .C(Cout[29]), .S(S[29])),
                       
                       tree30(.N(N30), .Cin(Cout29 ), .Cout(Cout30), .C(Cout[30]), .S(S[30])),
                       tree31(.N(N31), .Cin(Cout30 ), .Cout(Cout31), .C(Cout[31]), .S(S[31])),
                       tree32(.N(N32), .Cin(Cout31 ), .Cout(Cout32), .C(Cout[32]), .S(S[32])),
                       tree33(.N(N33), .Cin(Cout32 ), .Cout(Cout33), .C(Cout[33]), .S(S[33])),
                       tree34(.N(N34), .Cin(Cout33 ), .Cout(Cout34), .C(Cout[34]), .S(S[34])),
                       tree35(.N(N35), .Cin(Cout34 ), .Cout(Cout35), .C(Cout[35]), .S(S[35])),
                       tree36(.N(N36), .Cin(Cout35 ), .Cout(Cout36), .C(Cout[36]), .S(S[36])),
                       tree37(.N(N37), .Cin(Cout36 ), .Cout(Cout37), .C(Cout[37]), .S(S[37])),
                       tree38(.N(N38), .Cin(Cout37 ), .Cout(Cout38), .C(Cout[38]), .S(S[38])),
                       tree39(.N(N39), .Cin(Cout38 ), .Cout(Cout39), .C(Cout[39]), .S(S[39])),
                       
                       tree40(.N(N40), .Cin(Cout39 ), .Cout(Cout40), .C(Cout[40]), .S(S[40])),
                       tree41(.N(N41), .Cin(Cout40 ), .Cout(Cout41), .C(Cout[41]), .S(S[41])),
                       tree42(.N(N42), .Cin(Cout41 ), .Cout(Cout42), .C(Cout[42]), .S(S[42])),
                       tree43(.N(N43), .Cin(Cout42 ), .Cout(Cout43), .C(Cout[43]), .S(S[43])),
                       tree44(.N(N44), .Cin(Cout43 ), .Cout(Cout44), .C(Cout[44]), .S(S[44])),
                       tree45(.N(N45), .Cin(Cout44 ), .Cout(Cout45), .C(Cout[45]), .S(S[45])),
                       tree46(.N(N46), .Cin(Cout45 ), .Cout(Cout46), .C(Cout[46]), .S(S[46])),
                       tree47(.N(N47), .Cin(Cout46 ), .Cout(Cout47), .C(Cout[47]), .S(S[47])),
                       tree48(.N(N48), .Cin(Cout47 ), .Cout(Cout48), .C(Cout[48]), .S(S[48])),
                       tree49(.N(N49), .Cin(Cout48 ), .Cout(Cout49), .C(Cout[49]), .S(S[49])),                                              
                       
                       tree50(.N(N50), .Cin(Cout49 ), .Cout(Cout50), .C(Cout[50]), .S(S[50])),
                       tree51(.N(N51), .Cin(Cout50 ), .Cout(Cout51), .C(Cout[51]), .S(S[51])),
                       tree52(.N(N52), .Cin(Cout51 ), .Cout(Cout52), .C(Cout[52]), .S(S[52])),
                       tree53(.N(N53), .Cin(Cout52 ), .Cout(Cout53), .C(Cout[53]), .S(S[53])),
                       tree54(.N(N54), .Cin(Cout53 ), .Cout(Cout54), .C(Cout[54]), .S(S[54])),
                       tree55(.N(N55), .Cin(Cout54 ), .Cout(Cout55), .C(Cout[55]), .S(S[55])),
                       tree56(.N(N56), .Cin(Cout55 ), .Cout(Cout56), .C(Cout[56]), .S(S[56])),
                       tree57(.N(N57), .Cin(Cout56 ), .Cout(Cout57), .C(Cout[57]), .S(S[57])),
                       tree58(.N(N58), .Cin(Cout57 ), .Cout(Cout58), .C(Cout[58]), .S(S[58])),
                       tree59(.N(N59), .Cin(Cout58 ), .Cout(Cout59), .C(Cout[59]), .S(S[59])),   
                       
                       tree60(.N(N60), .Cin(Cout59 ), .Cout(Cout60), .C(Cout[60]), .S(S[60])),
                       tree61(.N(N61), .Cin(Cout60 ), .Cout(Cout61), .C(Cout[61]), .S(S[61])),
                       tree62(.N(N62), .Cin(Cout61 ), .Cout(Cout62), .C(Cout[62]), .S(S[62])),
                       tree63(.N(N63), .Cin(Cout62 ), .Cout(Cout63), .C(Cout[63]), .S(S[63]));
endmodule

module one_bit_Wallace_tree(
  input  [16:0] N,
  input  [13:0] Cin,

  output [13:0] Cout,
  output C,
  output S
);

  wire S00, S01, S02, S03, S04, S05, S06, S07, S08, S09, S10, S11, S12, S13;

  one_bit_full_adder adder00(.A(N[16]  ), .B(N[15]  ), .Cin(N[14]  ), .S(S00), .Cout(Cout[00])),
                     adder01(.A(N[13]  ), .B(N[12]  ), .Cin(N[11]  ), .S(S01), .Cout(Cout[01])),
                     adder02(.A(N[10]  ), .B(N[09]  ), .Cin(N[08]  ), .S(S02), .Cout(Cout[02])),
                     adder03(.A(N[07]  ), .B(N[06]  ), .Cin(N[05]  ), .S(S03), .Cout(Cout[03])),
                     adder04(.A(N[04]  ), .B(N[03]  ), .Cin(N[02]  ), .S(S04), .Cout(Cout[04])),
                     adder05(.A(S00    ), .B(S01    ), .Cin(S02    ), .S(S05), .Cout(Cout[05])),
                     adder06(.A(S03    ), .B(S04    ), .Cin(N[01]  ), .S(S06), .Cout(Cout[06])),
                     adder07(.A(N[00]  ), .B(Cin[00]), .Cin(Cin[01]), .S(S07), .Cout(Cout[07])),
                     adder08(.A(Cin[02]), .B(Cin[03]), .Cin(Cin[04]), .S(S08), .Cout(Cout[08])),
                     adder09(.A(S05    ), .B(S06    ), .Cin(S07    ), .S(S09), .Cout(Cout[09])),
                     adder10(.A(S08    ), .B(Cin[05]), .Cin(Cin[06]), .S(S10), .Cout(Cout[10])),
                     adder11(.A(S09    ), .B(S10    ), .Cin(Cin[07]), .S(S11), .Cout(Cout[11])),
                     adder12(.A(Cin[08]), .B(Cin[09]), .Cin(Cin[10]), .S(S12), .Cout(Cout[12])),
                     adder13(.A(S11    ), .B(S12    ), .Cin(Cin[11]), .S(S13), .Cout(Cout[13])),
                     adder14(.A(S13    ), .B(Cin[12]), .Cin(Cin[13]), .S(S  ), .Cout(C       ));
endmodule

module one_bit_full_adder(
  input A,
  input B,
  input Cin,
  
  output S,
  output Cout
);

  assign S = ~A & ~B & Cin | ~A & B & ~Cin | A & ~B & ~Cin | A & B & Cin;
  assign Cout = A & B |A & Cin | B & Cin;
 
endmodule

module final_adder(
  input  [63:0] A,
  input  [63:0] B,
  input  Cin,
  
  output [63:0] result
);


  assign result = A + B + Cin;
  
endmodule